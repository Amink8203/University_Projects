`timescale 1ns/1ns
module tb7();
    logic[14:0] t = 0;
    wire[3:0] out;
    ex7 CUT1(t,out);
    initial begin
      #200 t[0] = 1;
      #200 t[5] = 1;
      #200 t[1] = 1;
      #200 t[3] = 1;
      #200 t[2] = 1;
      #200 t[6] = 1;
      #200 t[4] = 1;
      #200 t[14] = 1;
      #200 t[8] = 1;
      #200 t[7] = 1;
      #200 t[12] = 1;
      #200 t[10] = 1;
      #200 t[11] = 1;
      #200 t[9] = 1;
      #200 t[13] = 1;

      #200 t[0] = 0;
      #200 t[5] = 0;
      #200 t[1] = 0;
      #200 t[3] = 0;
      #200 t[2] = 0;
      #200 t[6] = 0;
      #200 t[4] = 0;
      #200 t[14] = 0;
      #200 t[8] = 0;
      #200 t[7] = 0;
      #200 t[12] = 0;
      #200 t[10] = 0;
      #200 t[11] = 0;
      #200 t[9] = 0;
      #200 t[13] = 0;
      #250 $stop;
    end
endmodule



